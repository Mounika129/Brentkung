module a_bc_module(y,a,b,c);
input a,b,c;
output y;

assign y= a | ( b & c ) ;































endmodule 